* cir2
.options savecurrents

* Netlist

.include circuit2.txt

* Control Commands

.control
op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

echo  "op2_TAB"
print all
echo  "op2_END"

exit
.endc 
.end

