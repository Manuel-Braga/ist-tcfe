* T1
.options savecurrents

* Netlist

V0 1 0 0V
Va 2 1 5.06400320393
R1 2 3 1.00196314014
R2 3 4 2.082319235
R3 3 5 3.05798143645
R4 1 5 4.10496355098
R5 5 6 3.03658050119
R6 1 7 2.00356698935
R7 8 9 1.0495200477
Id 9 6 1.01960705059
VIc 7 8 0V
GIb 6 4 3 5 7.0260450587
HVc 5 9 VIc 8.35916956066


* Control Commands

.control
op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

echo  "op_TAB"
print all
echo  "op_END"


quit
.endc 

.end
